library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package bird_bitmap is
  type bird_rgb_pixel is array(0 to 2) of std_logic_vector(3 downto 0); -- [R,G,B]
  type bird_bitmap_type is array(0 to 19, 0 to 19) of bird_rgb_pixel;

  constant bird_bitmap : bird_bitmap_type := (
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("0001","0001","0001"), ("1111","1111","1111"), ("0100","0100","0100"), ("1111","1111","1111"), ("0111","0111","0111"), ("1111","1111","1111"), ("0010","0001","0001"), ("1111","1111","1111"), ("0001","0001","0001"), ("0000","0000","0000"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1011","0000"), ("1111","1011","0000"), ("0000","0000","0010"), ("0010","0010","0010"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1100","0000"), ("1111","1011","0000"), ("0010","0010","0010"), ("1111","1011","0000"), ("1111","1011","0000"), ("1110","1110","1110"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1100","0000"), ("1111","1011","0000"), ("1111","1100","0000"), ("0010","0010","0010"), ("1111","1011","0000"), ("1110","1110","1110"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1011","0000"), ("1111","1011","0000"), ("1111","1011","0000"), ("0010","0010","0010"), ("1111","1100","0000"), ("1111","1100","0000"), ("1110","0111","0000"), ("1110","0111","0000"), ("1110","0111","0000"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("0010","0010","0010"), ("1111","1010","0000"), ("0000","0000","0010"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"))
	);
end package bird_bitmap;