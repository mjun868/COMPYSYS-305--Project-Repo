constant bird_bitmap : bird_bitmap_type := (
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("0001","0001","0001"), ("1111","1111","1111"), ("0100","0100","0100"), ("1111","1111","1111"), ("0111","0111","0111"), ("1111","1111","1111"), ("0010","0001","0001"), ("1111","1111","1111"), ("0001","0001","0001"), ("0000","0000","0000"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1011","0000"), ("1111","1011","0000"), ("0000","0000","0010"), ("0010","0010","0010"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1100","0000"), ("1111","1011","0000"), ("0010","0010","0010"), ("1111","1011","0000"), ("1111","1011","0000"), ("1110","1110","1110"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1100","0000"), ("1111","1011","0000"), ("1111","1100","0000"), ("0010","0010","0010"), ("1111","1011","0000"), ("1110","1110","1110"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1011","0000"), ("1111","1011","0000"), ("1111","1011","0000"), ("0010","0010","0010"), ("1111","1100","0000"), ("1111","1100","0000"), ("1110","0111","0000"), ("1110","0111","0000"), ("1110","0111","0000"), ("1111","1111","1111"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("0010","0010","0010"), ("1111","1010","0000"), ("0000","0000","0010"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1010","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("0000","0000","0000"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111")),
    (("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"), ("1111","1111","1111"))
);