LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;



USE work.bird_bitmap.ALL;  -- Make sure you include your bird_bitmap package

ENTITY falling_bird IS
    PORT (
        clk, vert_sync        : IN std_logic;
        pixel_row, pixel_column : IN std_logic_vector(9 DOWNTO 0);
        red, green, blue        : OUT std_logic_vector(3 DOWNTO 0)
    );
END falling_bird;

ARCHITECTURE behavior OF falling_bird IS

  -- Sprite constants
  CONSTANT BIRD_X_POS  : integer := 80;         -- fixed horizontal position
  CONSTANT BIRD_WIDTH  : integer := 20;
  CONSTANT BIRD_HEIGHT : integer := 20;
  CONSTANT FALL_SPEED  : integer := 2;

  -- Signals for pixel control
  SIGNAL bird_on           : std_logic := '0';
  SIGNAL bird_y_pos        : integer := 200;
  SIGNAL pixel_x, pixel_y  : integer;
  SIGNAL bird_r, bird_g, bird_b : std_logic_vector(3 DOWNTO 0);

BEGIN

  -- Convert pixel_row and pixel_column to integers
  pixel_x <= to_integer(unsigned(pixel_column));
  pixel_y <= to_integer(unsigned(pixel_row));

  -- Sprite drawing logic
  PROCESS(clk)
    VARIABLE row_idx, col_idx : integer;
  BEGIN
    IF rising_edge(clk) THEN
      IF (pixel_x >= BIRD_X_POS AND pixel_x < BIRD_X_POS + BIRD_WIDTH) AND
         (pixel_y >= bird_y_pos AND pixel_y < bird_y_pos + BIRD_HEIGHT) THEN
         
        row_idx := pixel_y - bird_y_pos;
        col_idx := pixel_x - BIRD_X_POS;

        bird_on <= '1';

        bird_r <= bird_bitmap(row_idx, col_idx)(0);
        bird_g <= bird_bitmap(row_idx, col_idx)(1);
        bird_b <= bird_bitmap(row_idx, col_idx)(2);
      ELSE
        bird_on <= '0';
      END IF;
    END IF;
  END PROCESS;

  -- Gravity motion
  Move_Bird : PROCESS(vert_sync)
  BEGIN
    IF rising_edge(vert_sync) THEN
      IF bird_y_pos < (480 - BIRD_HEIGHT) THEN
        bird_y_pos <= bird_y_pos + FALL_SPEED;
      END IF;
    END IF;
  END PROCESS;

  -- RGB output (white background)
  red   <= bird_r WHEN bird_on = '1' ELSE "1111";
  green <= bird_g WHEN bird_on = '1' ELSE "1111";
  blue  <= bird_b WHEN bird_on = '1' ELSE "1111";

END behavior;

	
